LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE binary_instructions_package IS
    CONSTANT INSTR_WIDTH : NATURAL := 32;

    CONSTANT ADD_INSTR_RD : STD_LOGIC_VECTOR(5 - 1 DOWNTO 0) := B"00100";
    CONSTANT ADD_INSTR_RS1 : STD_LOGIC_VECTOR(5 - 1 DOWNTO 0) := B"00011";
    CONSTANT ADD_INSTR_RS2 : STD_LOGIC_VECTOR(5 - 1 DOWNTO 0) := B"00111";
    CONSTANT ADD_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"0000000" & ADD_INSTR_RS2 & ADD_INSTR_RS1 & B"000" & ADD_INSTR_RD & B"0110011"; -- d"10584627" -> R[rd] = R[rs1] + R[rs2] -> R[4] = R[3] + R[7]

    CONSTANT ADDI_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"00000000000000000000000000010011"; -- ADDI

    CONSTANT SLL_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"00000000000000000010000000110011"; -- SLL
    CONSTANT NOP_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"00000000000000000010000000010011"; -- ADDI
    CONSTANT LW_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"00000000000000000010000000000011"; -- LW
    CONSTANT BNE_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"00000000000000000001000000100011"; -- BNE
    CONSTANT BEQ_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"00000000000000000011000000100011"; -- BEQ
    CONSTANT SW_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"00000000000000000010000000100011"; -- SW
    CONSTANT J_INSTR_BINARY : STD_LOGIC_VECTOR(INSTR_WIDTH - 1 DOWNTO 0) := B"00000000000000000000000000000010"; -- J
END binary_instructions_package;
