LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE control_unit_outputs_package IS
    CONSTANT CONTROL_UNIT_OUTPUTS_WIDTH : NATURAL := 32;
    CONSTANT ADD_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000000100110"; -- X'2026, ADD
    CONSTANT SUB_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000001000110"; -- SUB
    CONSTANT SLL_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000010000110"; --  X'2086, SLL
    CONSTANT SRL_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000010100110"; -- SRL
    CONSTANT SLT_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000110000110"; -- SLT
    CONSTANT NOP_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000000000010"; -- NOP
    CONSTANT ADDI_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000001101110"; -- ADDI
    CONSTANT SLTI_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000110101110"; -- SLTI
    CONSTANT LB_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10001100001110"; -- LB
    CONSTANT LW_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10001011001110"; -- X'22CE, LW
    CONSTANT SB_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000100111010"; -- SB
    CONSTANT BNE_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10100101100010"; -- X'2962, BNE
    CONSTANT SW_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10000011111010"; -- X'20FA, SW
    CONSTANT BEQ_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"10010101000010"; -- X'2542, BEQ
    CONSTANT J_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"11110000000010"; -- X'3C02, J
    CONSTANT JAL_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"00110000000110"; -- JAL
    CONSTANT JARL_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"00110000001110"; -- JARL
    CONSTANT ECALL_CONTROL_UNIT_OUTPUT : STD_LOGIC_VECTOR(CONTROL_UNIT_OUTPUTS_WIDTH - 1 DOWNTO 0) := B"00000000000001"; -- ECALL
END control_unit_outputs_package;
